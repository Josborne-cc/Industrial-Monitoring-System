--Program: TDM_RECIEVER
--Purpose: Create TDM_RECIEVER
--Author: Josh Osborne 
--Date: November 16, 2014

--|Input Bit Stream of Data
--|Input
--|GPIO_0[1]
--|PIN_A13

--|Input Clock Pulse
--|CLK
--|24 MHz Clock
--|PIN_A12

--|HEX DISPLAYS
--|HEX3
--|HEX_3[0] |HEX_3[1] |HEX_3[2] |HEX_3[3] |HEX_3[4] |HEX_3[5] |HEX_3[6]
--|PIN_F4   |PIN_D5   |PIN_D6   |PIN_J4   |PIN_L8   |PIN_F3   |PIN_D4

--|HEX2
--|HEX_2[0] |HEX_2[1] |HEX_2[2] |HEX_2[3] |HEX_2[4] |HEX_2[5] |HEX_2[6]
--|PIN_G5   |PIN_G6   |PIN_C2   |PIN_C1   |PIN_E3   |PIN_E4   |PIN_D3

--|HEX1
--|HEX_1[0] |HEX_1[1] |HEX_1[2] |HEX_1[3] |HEX_1[4] |HEX_1[5] |HEX_1[6]
--|PIN_E1   |PIN_H6   |PIN_H5   |PIN_H4   |PIN_G3   |PIN_D2   |PIN_D1

--|HEX0
--|HEX_0[0] |HEX_0[1] |HEX_0[2] |HEX_0[3] |HEX_0[4] |HEX_0[5] |HEX_0[6]
--|PIN_J2   |PIN_J1   |PIN_H2   |PIN_H1   |PIN_F2   |PIN_F1   |PIN_E2

--|COUNT FOR OUPUT AS A DECREASING INTEGER
--| COUNT_ERROR_OUTPUT[7] | COUNT_ERROR_OUTPUT[6] | COUNT_ERROR_OUTPUT[5] | COUNT_ERROR_OUTPUT[4] | COUNT_ERROR_OUTPUT[3] | COUNT_ERROR_OUTPUT[2] | COUNT_ERROR_OUTPUT[1] | COUNT_ERROR_OUTPUT[0] |
--| LED_G7                | LED_G6                | LED_G5                | LED_G4                | LED_G3                | LED_RG2               | LED_G1                | LED_G0                |
--| PIN_Y21               | PIN_Y22               | PIN_W21               | PIN_W22               | PIN_V21               | PIN_V22               | PIN_U21               | PIN_U22               |

LIBRARY ieee;
	USE ieee.std_logic_1164.ALL;
	USE ieee.std_logic_unsigned.ALL;
	USE ieee.std_logic_ARITH.ALL;
	
 ENTITY TDM_RECIEVER IS
 
	PORT(CLK: IN STD_LOGIC;
		INPUT: IN STD_LOGIC;
		SYNC_CLK: IN STD_LOGIC;
		CONTROL: IN STD_LOGIC_VECTOR (1 	DOWNTO 0); --USED FOR HANDSHAKING WITH LARGE LCD DISPLAY
		DECODER_CLK: OUT STD_LOGIC;
		DISPLAY: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		HEX_0: OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
		HEX_1: OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
		HEX_2: OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
		HEX_3: OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
		OUTPUT_ERROR_COUNT: OUT STD_LOGIC_VECTOR (7 DOWNTO 0));
END TDM_RECIEVER;

ARCHITECTURE behaviour OF TDM_RECIEVER IS

	CONSTANT HIGH: STD_LOGIC := '1';
	CONSTANT LOW: STD_LOGIC := '0';
	CONSTANT VALUE_0: STD_LOGIC_VECTOR := "0000";
	CONSTANT VALUE_1: STD_LOGIC_VECTOR := "0001";
	CONSTANT VALUE_2: STD_LOGIC_VECTOR := "0010";
	CONSTANT VALUE_3: STD_LOGIC_VECTOR := "0011";
	CONSTANT VALUE_4: STD_LOGIC_VECTOR := "0100";
	CONSTANT VALUE_5: STD_LOGIC_VECTOR := "0101";
	CONSTANT VALUE_6: STD_LOGIC_VECTOR := "0110";
	CONSTANT VALUE_7: STD_LOGIC_VECTOR := "0111";
	CONSTANT VALUE_8: STD_LOGIC_VECTOR := "1000";
	CONSTANT VALUE_9: STD_LOGIC_VECTOR := "1001";
	CONSTANT VALUE_A: STD_LOGIC_VECTOR := "1010";
	CONSTANT VALUE_B: STD_LOGIC_VECTOR := "1011";
	CONSTANT VALUE_C: STD_LOGIC_VECTOR := "1100";
	CONSTANT VALUE_D: STD_LOGIC_VECTOR := "1101";
	CONSTANT VALUE_E: STD_LOGIC_VECTOR := "1110";
	CONSTANT VALUE_F: STD_LOGIC_VECTOR := "1111";
	CONSTANT HEX_DISPLAY_0: STD_LOGIC_VECTOR := "1000000";
	CONSTANT HEX_DISPLAY_1: STD_LOGIC_VECTOR := "1111001";
	CONSTANT HEX_DISPLAY_2: STD_LOGIC_VECTOR := "0100100";
	CONSTANT HEX_DISPLAY_3: STD_LOGIC_VECTOR := "0110000";
	CONSTANT HEX_DISPLAY_4: STD_LOGIC_VECTOR := "0011001";
	CONSTANT HEX_DISPLAY_5: STD_LOGIC_VECTOR := "0010010";
	CONSTANT HEX_DISPLAY_6: STD_LOGIC_VECTOR := "0000010";
	CONSTANT HEX_DISPLAY_7: STD_LOGIC_VECTOR := "1111000";
	CONSTANT HEX_DISPLAY_8: STD_LOGIC_VECTOR := "0000000";
	CONSTANT HEX_DISPLAY_9: STD_LOGIC_VECTOR := "0011000";
	CONSTANT HEX_DISPLAY_A: STD_LOGIC_VECTOR := "0001000";
	CONSTANT HEX_DISPLAY_B: STD_LOGIC_VECTOR := "0000011";
	CONSTANT HEX_DISPLAY_C: STD_LOGIC_VECTOR := "1000110";
	CONSTANT HEX_DISPLAY_D: STD_LOGIC_VECTOR := "0100001";
	CONSTANT HEX_DISPLAY_E: STD_LOGIC_VECTOR := "0000110";
	CONSTANT HEX_DISPLAY_F: STD_LOGIC_VECTOR := "0001110";
	CONSTANT HEX_DISPLAY_CLEAR: STD_LOGIC_VECTOR := "1111111";
	
	TYPE STATE IS (STATE0, STATE1, STATE2, STATE3, STATE4, STATE5, STATE6);
	SHARED VARIABLE PRESENTSTATE, NEXTSTATE: STATE;

	BEGIN
	
		PROCESS(SYNC_CLK)
			VARIABLE SYNC_CLK_COUNT: INTEGER := 0;
			VARIABLE SYNC_CLK_PULSE: STD_LOGIC := LOW;
			
			BEGIN
				IF  (RISING_EDGE(SYNC_CLK)) THEN
				
					SYNC_CLK_COUNT := SYNC_CLK_COUNT + 1;
					DECODER_CLK <= SYNC_CLK_PULSE;
					
					IF (SYNC_CLK_COUNT MOD 34 = 0) THEN
						SYNC_CLK_PULSE := SYNC_CLK_PULSE XOR HIGH;
					END IF;
					IF (SYNC_CLK_COUNT = 24000000) THEN
						SYNC_CLK_COUNT := 0;
					END IF;
				END IF;
			END PROCESS;
			
		PROCESS(CLK)
			VARIABLE TDM_VECTOR: STD_LOGIC_VECTOR (7 DOWNTO 0) := "00000000";
			VARIABLE TDM_VECTOR2: STD_LOGIC_VECTOR (7 DOWNTO 0) := "00000000";
			VARIABLE TDM_VECTOR3: STD_LOGIC_VECTOR (7 DOWNTO 0) := "00000000";
			VARIABLE SENSOR1_DATA: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
			VARIABLE SENSOR2_DATA: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
			VARIABLE TEMP: INTEGER := 0;
			VARIABLE ERROR_OUT: INTEGER := 0;
			VARIABLE DATA_COUNT: INTEGER := 0;
			VARIABLE ERROR_COUNT: INTEGER := 0;
			VARIABLE CORRECT_COUNT: INTEGER := 0;
			
			--Function to convert to HEX
			FUNCTION WRITEHEX(DATA: IN STD_LOGIC_VECTOR)
					RETURN STD_LOGIC_VECTOR IS
					VARIABLE VAR: STD_LOGIC_VECTOR(6 DOWNTO 0);
					
					BEGIN
						IF(DATA = VALUE_0) THEN
							VAR := HEX_DISPLAY_0;
						ELSIF(DATA = VALUE_1) THEN
							VAR := HEX_DISPLAY_1;
						ELSIF(DATA = VALUE_2) THEN
							VAR := HEX_DISPLAY_2;
						ELSIF(DATA = VALUE_3) THEN
							VAR := HEX_DISPLAY_3;
						ELSIF(DATA = VALUE_4) THEN
							VAR := HEX_DISPLAY_4;
						ELSIF(DATA = VALUE_5) THEN
							VAR := HEX_DISPLAY_5;
						ELSIF(DATA = VALUE_6) THEN
							VAR := HEX_DISPLAY_6;
						ELSIF(DATA = VALUE_7) THEN
							VAR := HEX_DISPLAY_7;
						ELSIF(DATA = VALUE_8) THEN
							VAR := HEX_DISPLAY_8;
						ELSIF(DATA = VALUE_9) THEN
							VAR := HEX_DISPLAY_9;
						ELSIF(DATA = VALUE_A) THEN
							VAR := HEX_DISPLAY_A;
						ELSIF(DATA = VALUE_B) THEN
							VAR := HEX_DISPLAY_B;
						ELSIF(DATA = VALUE_C) THEN
							VAR := HEX_DISPLAY_C;
						ELSIF(DATA = VALUE_D) THEN
							VAR := HEX_DISPLAY_D;
						ELSIF(DATA = VALUE_E) THEN
							VAR := HEX_DISPLAY_E;
						ELSIF(DATA = VALUE_F) THEN
							VAR := HEX_DISPLAY_F;
						END IF;
						
						RETURN VAR;
					END WRITEHEX;
			
			BEGIN 

				IF (RISING_EDGE (CLK)) THEN
				--Goes to the next state
				PRESENTSTATE := NEXTSTATE; 
				
				CASE PRESENTSTATE IS
				
					WHEN STATE0 =>
						--Collect Data
						TDM_VECTOR(7 DOWNTO 1) := TDM_VECTOR (6 DOWNTO 0); --Move the input on bit to the left
						TDM_VECTOR(0) := INPUT; --Saves the last input for these 8 bits
						
						TEMP := (ERROR_COUNT /  CORRECT_COUNT) * 100;
						ERROR_OUT := TEMP;
						
						--Converts the integer into a vector
						OUTPUT_ERROR_COUNT <= "00000000";
						--OUTPUT_ERROR_COUNT <= CONV_STD_LOGIC_VECTOR(TEMP, 8);
						
						IF (TDM_VECTOR = x"FF") THEN	
							TDM_VECTOR (7 DOWNTO 0) := "00000000";
							--Sync frame is found 
							NEXTSTATE := STATE1;
						ELSE
							NEXTSTATE := STATE0;
						END IF;
						
					WHEN STATE1 =>
						--Gets the second 0xFF data from sender
						DATA_COUNT := DATA_COUNT + 1;
						IF (DATA_COUNT < 9) THEN
							TDM_VECTOR(7 DOWNTO 1) := TDM_VECTOR(6 DOWNTO 0);
							TDM_VECTOR(0) := INPUT;
							NEXTSTATE := STATE1;
						END IF;
						
						IF (DATA_COUNT = 8) THEN
							DATA_COUNT := 0;
							
							IF (TDM_VECTOR = x"FF") THEN
								TDM_VECTOR (7 DOWNTO 0) := "00000000";
								NEXTSTATE := STATE2;
							ELSIF (TDM_VECTOR /= x"FF") THEN
								TDM_VECTOR (7 DOWNTO 0) := "00000000";
								NEXTSTATE := STATE0;
							END IF;
							
						END IF;
							
					WHEN STATE2 =>
						--Gets Sensor 1 data
						DATA_COUNT := DATA_COUNT + 1;
						
						--Collect 16-bits of data
						IF (DATA_COUNT <= 8) THEN
							TDM_VECTOR(7 DOWNTO 1) := TDM_VECTOR(6 DOWNTO 0);
							TDM_VECTOR(0) := INPUT;
							NEXTSTATE := STATE2;
						ELSIF (DATA_COUNT >= 9) THEN
							TDM_VECTOR2(7 DOWNTO 1) := TDM_VECTOR2(6 DOWNTO 0);
							TDM_VECTOR2(0) := INPUT;
							NEXTSTATE := STATE2;
						END IF;
						
						IF (DATA_COUNT = 16) THEN
							DATA_COUNT := 0;
							--XOR the 16bits we need to get 0xFF
							TDM_VECTOR3 := TDM_VECTOR XOR TDM_VECTOR2;
							
							IF(TDM_VECTOR3 = x"FF") THEN
								CORRECT_COUNT := CORRECT_COUNT + 1;
								SENSOR1_DATA := TDM_VECTOR;
								HEX_2 <= WRITEHEX(TDM_VECTOR(3 DOWNTO 0));
								HEX_3 <= WRITEHEX(TDM_VECTOR(7 DOWNTO 4));
								TDM_VECTOR (7 DOWNTO 0) := "00000000";
								NEXTSTATE := STATE3;
							ELSE
								ERROR_COUNT := ERROR_COUNT + 1;
								TDM_VECTOR (7 DOWNTO 0) := "00000000";
								NEXTSTATE := STATE3;
							END IF;
						END IF;
						
					WHEN STATE3 =>
							--Gets 0xAA
							DATA_COUNT := DATA_COUNT + 1;
							
							IF (DATA_COUNT < 9) THEN
								TDM_VECTOR(7 DOWNTO 1) := TDM_VECTOR(6 DOWNTO 0);
								TDM_VECTOR(0) := INPUT;
								NEXTSTATE := STATE3;
							END IF;
							
							IF (DATA_COUNT = 8) THEN
								DATA_COUNT := 0;
								
								IF (TDM_VECTOR = x"AA") THEN
									TDM_VECTOR (7 DOWNTO 0) := "00000000";
									NEXTSTATE := STATE4;
								ELSE
									TDM_VECTOR (7 DOWNTO 0) := "00000000";
									NEXTSTATE := STATE0;
								END IF;
							END IF;
							
					WHEN STATE4 =>
						--Gets Sensor 2 data
						DATA_COUNT := DATA_COUNT + 1;
						
						IF (DATA_COUNT <= 8) THEN
							TDM_VECTOR(7 DOWNTO 1) := TDM_VECTOR(6 DOWNTO 0);
							TDM_VECTOR(0) := INPUT;
							NEXTSTATE := STATE4;
						ELSIF (DATA_COUNT >= 9) THEN
							TDM_VECTOR2(7 DOWNTO 1) := TDM_VECTOR2(6 DOWNTO 0);
							TDM_VECTOR2(0) := INPUT;
							NEXTSTATE := STATE4;
						END IF;
							
						IF (DATA_COUNT = 16) THEN
							DATA_COUNT := 0;
							
							TDM_VECTOR3 := TDM_VECTOR XOR TDM_VECTOR2;
							
							IF(TDM_VECTOR3 = x"FF") THEN
								CORRECT_COUNT := CORRECT_COUNT + 1;
								SENSOR2_DATA := TDM_VECTOR;
								HEX_0 <= WRITEHEX(TDM_VECTOR(3 DOWNTO 0));
								HEX_1 <= WRITEHEX(TDM_VECTOR(7 DOWNTO 4));
								TDM_VECTOR (7 DOWNTO 0) := "00000000";
								NEXTSTATE := STATE5;
							ELSE
								ERROR_COUNT := ERROR_COUNT + 1;
								TDM_VECTOR (7 DOWNTO 0) := "00000000";
								NEXTSTATE := STATE5;
							END IF;
						END IF;
						
					WHEN STATE5 =>
							
							DATA_COUNT := DATA_COUNT + 1;
							--Gets 0xAA
							IF (DATA_COUNT < 9) THEN
								TDM_VECTOR(7 DOWNTO 1) := TDM_VECTOR(6 DOWNTO 0);
								TDM_VECTOR(0) := INPUT;
								NEXTSTATE := STATE5;
							END IF;
							
							IF (DATA_COUNT = 8) THEN
								DATA_COUNT := 0;
								
								IF (TDM_VECTOR = x"AA") THEN
									TDM_VECTOR (7 DOWNTO 0) := "00000000";
									--NEXTSTATE := STATE0;
									NEXTSTATE := STATE6;
								ELSE
									TDM_VECTOR (7 DOWNTO 0) := "00000000";
									NEXTSTATE := STATE0;
								END IF;
							END IF;
					
					--HANDSHAKING WITH LCD DISPLAY
					WHEN STATE6 =>
						IF (CONTROL = "00") THEN
							DISPLAY <= "11111111";
							NEXTSTATE := STATE0;
						ELSIF (CONTROL = "01") THEN
							DISPLAY <= SENSOR1_DATA;
							NEXTSTATE := STATE6;
						ELSIF(CONTROL = "10") THEN
							DISPLAY <= SENSOR2_DATA;
							NEXTSTATE := STATE6;
						ELSIF(CONTROL = "11") THEN
							--DISPLAY <= CONV_STD_LOGIC_VECTOR(ERROR_OUT, 8);
							DISPLAY <= "00000000";
							NEXTSTATE := STATE6;
						END IF;
					
				END CASE;
				END IF;
		END PROCESS;
	END;

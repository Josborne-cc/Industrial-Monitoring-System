--Program: Time Division Multiplexer
--Purpose: Sender For Project
--Author: Josh Osborne, William Veldhuis and Colin Stanley
--Date: September 25, 2014


--|Main Clock Pulse
--|CLK
--|24 MHz Clock
--|PIN_A12

--|Sensor 1 Data Input
--|INPUT_SENSOR1[0] |INPUT_SENSOR1[1] |INPUT_SENSOR1[2] |INPUT_SENSOR1[3] |INPUT_SENSOR1[4] |INPUT_SENSOR1[5] |INPUT_SENSOR1[6] |INPUT_SENSOR1[7]
--|GPIO_0[11]       |GPIO_0[13]       |GPIO_0[15]       |GPIO_0[17]       |GPIO_0[19]       |GPIO_0[21]       |GPIO_0[23]       |GPIO_0[25]        
--|PIN_B18          |PIN_B19          |PIN_B20          |PIN_C22          |PIN_D22          |PIN_E22          |PIN_F22          |PIN_G22          

--|Sensor 2 Data Input
--|INPUT_SENSOR2[0] |INPUT_SENSOR2[1] |INPUT_SENSOR2[2] |INPUT_SENSOR2[3] |INPUT_SENSOR2[4] |INPUT_SENSOR2[5] |INPUT_SENSOR2[6] |INPUT_SENSOR2[7]
--|GPIO_0[10]       |GPIO_0[12]       |GPIO_0[14]       |GPIO_0[16]       |GPIO_0[18]       |GPIO_0[20]       |GPIO_0[22]       |GPIO_0[24]        
--|PIN_A18          |PIN_A19          |PIN_A20          |PIN_C21          |PIN_D21          |PIN_E21          |PIN_F21          |PIN_G21          

--|HEX DISPLAYS
--|HEX3
--|HEX_3[0] |HEX_3[1] |HEX_3[2] |HEX_3[3] |HEX_3[4] |HEX_3[5] |HEX_3[6]
--|PIN_F4   |PIN_D5   |PIN_D6   |PIN_J4   |PIN_L8   |PIN_F3   |PIN_D4

--|HEX2
--|HEX_2[0] |HEX_2[1] |HEX_2[2] |HEX_2[3] |HEX_2[4] |HEX_2[5] |HEX_2[6]
--|PIN_G5   |PIN_G6   |PIN_C2   |PIN_C1   |PIN_E3   |PIN_E4   |PIN_D3

--|HEX1
--|HEX_1[0] |HEX_1[1] |HEX_1[2] |HEX_1[3] |HEX_1[4] |HEX_1[5] |HEX_1[6]
--|PIN_E1   |PIN_H6   |PIN_H5   |PIN_H4   |PIN_G3   |PIN_D2   |PIN_D1

--|HEX0
--|HEX_0[0] |HEX_0[1] |HEX_0[2] |HEX_0[3] |HEX_0[4] |HEX_0[5] |HEX_0[6]
--|PIN_J2   |PIN_J1   |PIN_H2   |PIN_H1   |PIN_F2   |PIN_F1   |PIN_E2

--|Ouput Bit Stream of Data
--|OUPUT_DATA
--|GPIO_0[1]
--|PIN_A13

--|Output Clock Pulse
--|CLK_PULSE_OUT
--|GPIO_0[6]
--|PIN_A16



LIBRARY ieee;
	USE ieee.std_logic_1164.ALL;
	
ENTITY TDM_SENDER IS

	PORT (CLK: IN STD_LOGIC;
			INPUT_SENSOR1: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
			INPUT_SENSOR2: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
			HEX_0: OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
			HEX_1: OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
			HEX_2: OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
			HEX_3: OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
			CLK_PULSE_OUT: OUT STD_LOGIC;
			OUTPUT_DATA : OUT STD_LOGIC);
END TDM_SENDER;

ARCHITECTURE behaviour OF TDM_SENDER IS

	CONSTANT HIGH: STD_LOGIC := '1';
	CONSTANT LOW: STD_LOGIC := '0';
	CONSTANT VALUE_0: STD_LOGIC_VECTOR := "0000";
	CONSTANT VALUE_1: STD_LOGIC_VECTOR := "0001";
	CONSTANT VALUE_2: STD_LOGIC_VECTOR := "0010";
	CONSTANT VALUE_3: STD_LOGIC_VECTOR := "0011";
	CONSTANT VALUE_4: STD_LOGIC_VECTOR := "0100";
	CONSTANT VALUE_5: STD_LOGIC_VECTOR := "0101";
	CONSTANT VALUE_6: STD_LOGIC_VECTOR := "0110";
	CONSTANT VALUE_7: STD_LOGIC_VECTOR := "0111";
	CONSTANT VALUE_8: STD_LOGIC_VECTOR := "1000";
	CONSTANT VALUE_9: STD_LOGIC_VECTOR := "1001";
	CONSTANT VALUE_A: STD_LOGIC_VECTOR := "1010";
	CONSTANT VALUE_B: STD_LOGIC_VECTOR := "1011";
	CONSTANT VALUE_C: STD_LOGIC_VECTOR := "1100";
	CONSTANT VALUE_D: STD_LOGIC_VECTOR := "1101";
	CONSTANT VALUE_E: STD_LOGIC_VECTOR := "1110";
	CONSTANT VALUE_F: STD_LOGIC_VECTOR := "1111";
	CONSTANT HEX_DISPLAY_0: STD_LOGIC_VECTOR := "1000000";
	CONSTANT HEX_DISPLAY_1: STD_LOGIC_VECTOR := "1111001";
	CONSTANT HEX_DISPLAY_2: STD_LOGIC_VECTOR := "0100100";
	CONSTANT HEX_DISPLAY_3: STD_LOGIC_VECTOR := "0110000";
	CONSTANT HEX_DISPLAY_4: STD_LOGIC_VECTOR := "0011001";
	CONSTANT HEX_DISPLAY_5: STD_LOGIC_VECTOR := "0010010";
	CONSTANT HEX_DISPLAY_6: STD_LOGIC_VECTOR := "0000010";
	CONSTANT HEX_DISPLAY_7: STD_LOGIC_VECTOR := "1111000";
	CONSTANT HEX_DISPLAY_8: STD_LOGIC_VECTOR := "0000000";
	CONSTANT HEX_DISPLAY_9: STD_LOGIC_VECTOR := "0011000";
	CONSTANT HEX_DISPLAY_A: STD_LOGIC_VECTOR := "0001000";
	CONSTANT HEX_DISPLAY_B: STD_LOGIC_VECTOR := "0000011";
	CONSTANT HEX_DISPLAY_C: STD_LOGIC_VECTOR := "1000110";
	CONSTANT HEX_DISPLAY_D: STD_LOGIC_VECTOR := "0100001";
	CONSTANT HEX_DISPLAY_E: STD_LOGIC_VECTOR := "0000110";
	CONSTANT HEX_DISPLAY_F: STD_LOGIC_VECTOR := "0001110";
	CONSTANT HEX_DISPLAY_CLEAR: STD_LOGIC_VECTOR := "1111111";
	CONSTANT MAX: STD_LOGIC_VECTOR (7 DOWNTO 0) := x"FE";
	CONSTANT MIN: STD_LOGIC_VECTOR (7 DOWNTO 0) := x"01";
	CONSTANT SYNCH_BIT1: STD_LOGIC_VECTOR (7 DOWNTO 0) := x"FF";
	CONSTANT SYNCH_BIT2: STD_LOGIC_VECTOR (7 DOWNTO 0) := x"AA";
	TYPE STATE IS (STATE0, STATE1, STATE2, STATE3, STATE4, STATE5, STATE6, STATE7);
	SIGNAL PRESENTSTATE, NEXTSTATE: STATE;
	SHARED VARIABLE TDM_FRAME: STD_LOGIC_VECTOR (63 DOWNTO 0);
	
	BEGIN

	PROCESS(CLK)
	
		VARIABLE CLK_COUNT: INTEGER := 0;
		VARIABLE CLK_PULSE: STD_LOGIC := '0';
		VARIABLE ELEMENT: INTEGER := 64;
		BEGIN
			IF (RISING_EDGE(CLK)) THEN
			
				CLK_COUNT := CLK_COUNT + 1;
				CLK_PULSE_OUT <= CLK_PULSE;	--Sends the clock pulse to the reciever
					
				IF (CLK_COUNT MOD  16 = 0) THEN
					CLK_PULSE := CLK_PULSE XOR '1'; --Create a pulse which the reciever can sink to
				END IF;
				
				IF (CLK_COUNT = 1000) THEN
						PRESENTSTATE <= NEXTSTATE;
						OUTPUT_DATA <= TDM_FRAME(ELEMENT); --Sends the sensor information
						ELEMENT := ELEMENT - 1;
						CLK_COUNT := 0;
						IF (ELEMENT = 0) THEN
							ELEMENT := 64;
						END IF;
						
					END IF;
				
				
			END IF;
	END PROCESS;
	
		PROCESS (PRESENTSTATE, INPUT_SENSOR1, INPUT_SENSOR2)
		
			VARIABLE NORMAL_DATA_SENSOR1: STD_LOGIC_VECTOR (7 DOWNTO 0);
			VARIABLE NORMAL_DATA_SENSOR2: STD_LOGIC_VECTOR (7 DOWNTO 0);
			VARIABLE INVERTED_DATA_SENSOR1: STD_LOGIC_VECTOR (7 DOWNTO 0);
			VARIABLE INVERTED_DATA_SENSOR2: STD_LOGIC_VECTOR (7 DOWNTO 0);

				--FUNCTION ALLOWS FOR WRITING TO HEX DISPLAYS
				FUNCTION WRITEHEX(DATA: IN STD_LOGIC_VECTOR)
					RETURN STD_LOGIC_VECTOR IS
					VARIABLE VAR: STD_LOGIC_VECTOR(6 DOWNTO 0);
					
					BEGIN
						IF(DATA = VALUE_0) THEN
							VAR := HEX_DISPLAY_0;
						ELSIF(DATA = VALUE_1) THEN
							VAR := HEX_DISPLAY_1;
						ELSIF(DATA = VALUE_2) THEN
							VAR := HEX_DISPLAY_2;
						ELSIF(DATA = VALUE_3) THEN
							VAR := HEX_DISPLAY_3;
						ELSIF(DATA = VALUE_4) THEN
							VAR := HEX_DISPLAY_4;
						ELSIF(DATA = VALUE_5) THEN
							VAR := HEX_DISPLAY_5;
						ELSIF(DATA = VALUE_6) THEN
							VAR := HEX_DISPLAY_6;
						ELSIF(DATA = VALUE_7) THEN
							VAR := HEX_DISPLAY_7;
						ELSIF(DATA = VALUE_8) THEN
							VAR := HEX_DISPLAY_8;
						ELSIF(DATA = VALUE_9) THEN
							VAR := HEX_DISPLAY_9;
						ELSIF(DATA = VALUE_A) THEN
							VAR := HEX_DISPLAY_A;
						ELSIF(DATA = VALUE_B) THEN
							VAR := HEX_DISPLAY_B;
						ELSIF(DATA = VALUE_C) THEN
							VAR := HEX_DISPLAY_C;
						ELSIF(DATA = VALUE_D) THEN
							VAR := HEX_DISPLAY_D;
						ELSIF(DATA = VALUE_E) THEN
							VAR := HEX_DISPLAY_E;
						ELSIF(DATA = VALUE_F) THEN
							VAR := HEX_DISPLAY_F;
						END IF;
						
						RETURN VAR;
					END WRITEHEX;
			
			BEGIN 
			 
				
					CASE PRESENTSTATE IS
					
						WHEN STATE0 => 
								--Places 0xFF in the vector
								TDM_FRAME (63 DOWNTO 56) := SYNCH_BIT1; 
							
							NEXTSTATE <= STATE1;
							
						WHEN STATE1 => 
								--Places 0xFF in the vector for the second time
								TDM_FRAME (55 DOWNTO 48) := SYNCH_BIT1;

							NEXTSTATE <= STATE2;
							
						WHEN STATE2 =>
							--RESTRICTS INPUT FROM EVER BEING FF OR 00
							IF (INPUT_SENSOR1 = x"FF") THEN
								NORMAL_DATA_SENSOR1 := MAX;
								INVERTED_DATA_SENSOR1 := MIN;
							ELSIF (INPUT_SENSOR1 = x"00") THEN
								NORMAL_DATA_SENSOR1 := MIN;
								INVERTED_DATA_SENSOR1 := MAX;
							ELSE
								NORMAL_DATA_SENSOR1 := INPUT_SENSOR1;
								INVERTED_DATA_SENSOR1 := NOT(INPUT_SENSOR1);
							END IF;
							
							HEX_2 <= WRITEHEX(NORMAL_DATA_SENSOR1(3 DOWNTO 0));
							HEX_3 <= WRITEHEX(NORMAL_DATA_SENSOR1(7 DOWNTO 4));
							
							--Places the data from sensor 1 into the vector
							--FOR I IN 7 DOWNTO 0 LOOP
								TDM_FRAME(47 DOWNTO 40) := NORMAL_DATA_SENSOR1;
							--END LOOP;
							
							NEXTSTATE <= STATE3;
							
						WHEN STATE3 =>
								--Places the inverting data into the vector
								TDM_FRAME (39 DOWNTO 32) := INVERTED_DATA_SENSOR1;
			
							NEXTSTATE <= STATE4;
							
						WHEN STATE4 => 
							--Places 0xAA
							TDM_FRAME (31 DOWNTO 24) := SYNCH_BIT2;
							
							NEXTSTATE <= STATE5;
							
						WHEN STATE5 =>
							--RESTRICTS INPUT FROM EVER BEING FF OR 00
							IF (INPUT_SENSOR2 = x"FF") THEN
								NORMAL_DATA_SENSOR2 := x"FE";
								INVERTED_DATA_SENSOR2 := x"01";
							ELSIF (INPUT_SENSOR2 = x"00") THEN
								NORMAL_DATA_SENSOR2 := x"01";
								INVERTED_DATA_SENSOR2 := x"FE";
							ELSE
								NORMAL_DATA_SENSOR2 := INPUT_SENSOR2;
								INVERTED_DATA_SENSOR2 := NOT(INPUT_SENSOR2);
							END IF;
							
							HEX_0 <= WRITEHEX(NORMAL_DATA_SENSOR2(3 DOWNTO 0));
							HEX_1 <= WRITEHEX(NORMAL_DATA_SENSOR2(7 DOWNTO 4));
							--Places the data from sensor 2 into the vector
							TDM_FRAME (23 DOWNTO 16) := NORMAL_DATA_SENSOR2;
							
							NEXTSTATE <= STATE6;
							
						WHEN STATE6 => 
							--Places the inverting data into the vector
							TDM_FRAME (15 DOWNTO 8) := INVERTED_DATA_SENSOR2;
						
							NEXTSTATE <= STATE7;
							
						WHEN STATE7 => 
							--Places 0xAA after the second sensor data
							TDM_FRAME (7 DOWNTO 0) := SYNCH_BIT2;
							
							NEXTSTATE <= STATE0;
							
					END CASE;
			END PROCESS;
		END;
